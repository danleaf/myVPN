//x32+x26+x23+x22+x16+x12+x11+x10+x8+x7+x5+x4+x2+x1+1

module crc
#(parameter INIT = 32'hFFFFFFFF)
(
	input clk,rst_n,en,
	input [7:0] d,
	output [31:0] crc
);
	reg [31:0] r;
	wire sig;
	
	assign crc = r;
	
	initial
	begin
		r = INIT;
	end	
	
	always@(posedge clk or negedge rst_n)
	if(!rst_n)
		r <= INIT;
	else if(en)
	begin
		r[31] <= r[23] ^ r[29] ^ d[2];
		r[30] <= r[22] ^ r[28] ^ r[31] ^ d[0] ^ d[3];
		r[29] <= r[21] ^ r[27] ^ r[30] ^ r[31] ^ d[0] ^ d[1] ^ d[4];
		r[28] <= r[20] ^ r[30] ^ r[29] ^ r[26] ^ d[1] ^ d[2] ^ d[5];
		r[27] <= r[19] ^ r[25] ^ r[28] ^ r[29] ^ r[31] ^ d[0] ^ d[2] ^ d[3] ^ d[6];
		r[26] <= r[18] ^ r[24] ^ r[27] ^ r[28] ^ r[30] ^ d[1] ^ d[3] ^ d[4] ^ d[7];
		r[25] <= r[17] ^ r[26] ^ r[27] ^ d[4] ^ d[5];
		r[24] <= r[16] ^ r[25] ^ r[26] ^ r[31] ^ d[0] ^ d[5] ^ d[6];
		
		r[23] <= r[15] ^ r[24] ^ r[25] ^ r[30] ^ d[1] ^ d[6] ^ d[7];
		r[22] <= r[14] ^ r[24] ^ d[7];
		r[21] <= r[13] ^ r[29] ^ d[2];
		r[20] <= r[12] ^ r[28] ^ d[3];
		r[19] <= r[11] ^ r[27] ^ r[31] ^ d[0] ^ d[4];
		r[18] <= r[10] ^ r[26] ^ r[30] ^ r[31] ^ d[0] ^ d[1] ^ d[5];
		r[17] <= r[9] ^ r[25] ^ r[29] ^ r[30] ^ d[1] ^ d[2] ^ d[6];
		r[16] <= r[8] ^ r[24] ^ r[28] ^ r[29] ^ d[2] ^ d[3] ^ d[7];
		
		r[15] <= r[7] ^ r[27] ^ r[28] ^ r[29] ^ r[31] ^ d[0] ^ d[2] ^ d[3] ^ d[4];
		r[14] <= r[6] ^ r[26] ^ r[27] ^ r[28] ^ r[30] ^ r[31] ^ d[0] ^ d[1] ^ d[3] ^ d[4] ^ d[5];
		r[13] <= r[5] ^ r[25] ^ r[26] ^ r[27] ^ r[29] ^ r[30] ^ r[31] ^ d[0] ^ d[1] ^ d[2] ^ d[4] ^ d[5] ^ d[6];
		r[12] <= r[4] ^ r[24] ^ r[25] ^ r[26] ^ r[28] ^ r[29] ^ r[30] ^ d[1] ^ d[2] ^ d[3] ^ d[5] ^ d[6] ^ d[7];
		r[11] <= r[3] ^ r[24] ^ r[25] ^ r[27] ^ r[28] ^ d[3] ^ d[4] ^ d[6] ^ d[7];
		r[10] <= r[2] ^ r[24] ^ r[26] ^ r[27] ^ r[29] ^ d[2] ^ d[4] ^ d[5] ^ d[7];
		r[9] <= r[1] ^ r[25] ^ r[26] ^ r[28] ^ r[29] ^ d[2] ^ d[3] ^ d[5] ^ d[6];
		r[8] <= r[0] ^ r[24] ^ r[25] ^ r[27] ^ r[28] ^ d[3] ^ d[4] ^ d[6] ^ d[7];
		
		r[7] <= r[24] ^ r[26] ^ r[27] ^ r[29] ^ r[31] ^ d[0] ^ d[2] ^ d[4] ^ d[5] ^ d[7];
		r[6] <= r[25] ^ r[26] ^ r[28] ^ r[29] ^ r[30] ^ r[31] ^ d[0] ^ d[1] ^ d[2] ^ d[3] ^ d[5] ^ d[6];
		r[5] <= r[24] ^ r[25] ^ r[27] ^ r[28] ^ r[29] ^ r[30] ^ r[31] ^ d[0] ^ d[1] ^ d[2] ^ d[3] ^ d[4] ^ d[6] ^ d[7];
		r[4] <= r[24] ^ r[26] ^ r[27] ^ r[28] ^ r[30] ^ d[1] ^ d[3] ^ d[4] ^ d[5] ^ d[7];
		r[3] <= r[25] ^ r[26] ^ r[27] ^ r[31] ^ d[0] ^ d[4] ^ d[5] ^ d[6];
		r[2] <= r[24] ^ r[25] ^ r[26] ^ r[30] ^ r[31] ^ d[0] ^ d[1] ^ d[5] ^ d[6] ^ d[7];
		r[1] <= r[24] ^ r[25] ^ r[30] ^ r[31] ^ d[0] ^ d[1] ^ d[6] ^ d[7];
		r[0] <= r[24] ^ r[30] ^ d[1] ^ d[7];
	end

endmodule
